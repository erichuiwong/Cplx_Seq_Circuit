`include "dff.v"
module 8bitreg (
	//calls the 1 bit flip flop 8 times
);


